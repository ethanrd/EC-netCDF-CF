netcdf corridor_volume {
  dimensions:
      time = UNLIMITED ; // currently 11
      vol_width = 3 ;
      lat = 3 ;
      lon = 4 ;
      level = 5 ;
  variables:
      int time(time) ;
          time:units = "minutes since 2018-03-12T09:00Z"
      double lat(time, level, lat, lon, vol_width) ;
          lat:units = "degrees_north" ;
          lat:standard_name = "latitude" ;
      double lon(time, level, lat, lon, vol_width) ;
          lat:units = "degrees_east" ;
          lat:standard_name = "longitude" ;
      double level(time, level, lat, lon, vol_width) ;
          level:units = "meters" ;
          level:standard_name = "" ;
      double temp(time, level, lat, lon, vol_width) ;
          temp:units = "degC" ;
          temp:standard_name = "temperature" ;
//  data:
//      time = 0, 30, 60, 90, 120, 150, 180, 210, 240, 270, 300 ;
//      lat =
}