netcdf corridor_volume_separate {
  dimensions:
      time = UNLIMITED ; // currently 11
      vol_width = 3 ;
      vol_lat = 3 ;
      vol_lon = 4 ;
      vol_level = 5 ;
  variables:
      int time(time) ;
          time:units = "minutes since 2018-03-12T09:00Z"
      double traj_lat(time) ;
          traj_lat:units = "degrees_north" ;
          traj_lat:standard_name = "latitude" ;
      double traj_lon(time) ;
          traj_lat:units = "degrees_east" ;
          traj_lat:standard_name = "longitude" ;
      double traj_level(time) ;
          traj_level:units = "meters" ;
          traj_level:standard_name = "" ;


      double vol_lat(time, vol_level, vol_lat, vol_lon, vol_width) ;
          lat:units = "degrees_north" ;
          lat:standard_name = "latitude" ;
      double vol_lon(time, vol_level, vol_lat, vol_lon, vol_width) ;
          lat:units = "degrees_east" ;
          lat:standard_name = "longitude" ;
      double vol_level(time, vol_level, vol_lat, vol_lon, vol_width) ;
          level:units = "meters" ;
          level:standard_name = "" ;
      double temp(time, vol_level, vol_lat, vol_lon, vol_width) ;
          temp:units = "degC" ;
          temp:standard_name = "temperature" ;
//  data:
//      time = 0, 30, 60, 90, 120, 150, 180, 210, 240, 270, 300 ;
//      lat =
}
netcdf corridor_volume_separate {
  dimensions:
      time = UNLIMITED ; // currently 11
      lat = 3 ;
      lon = 4 ;
      level = 5 ;
  variables:
      int time(time) ;
          time:units = "minutes since 2018-03-12T09:00Z"
      double lat(time, level, lat, lon) ;
          lat:units = "degrees_north" ;
          lat:standard_name = "latitude" ;
      double lon(time, level, lat, lon) ;
          lat:units = "degrees_east" ;
          lat:standard_name = "longitude" ;
      double level(time, level, lat, lon) ;
          level:units = "meters" ;
          level:standard_name = "" ;
      double temp(time, level, lat, lon) ;
          temp:units = "degC" ;
          temp:standard_name = "temperature" ;
//  data:
//      time = 0, 30, 60, 90, 120, 150, 180, 210, 240, 270, 300 ;
//      lat =
}